output wire_out;

and a1(wire_out, , );
or o1(wire_out, , );
endmodule //\Users\epics\Documents\GitHub\uiverilog\output.v
