output ;

and a1(, , );
or o1(, , );
endmodule //\Users\epics\Documents\GitHub\uiverilog\output.v
